module top;
	initial begin
			$display("Practicing the version control");
			$display("Amend");
		$display("Going to pull");
	end
endmodule
