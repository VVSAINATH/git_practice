module top;
	initial begin
			$display("Practicing the version control");
			$display("Amend");
	end
endmodule
