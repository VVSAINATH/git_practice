module top;
	initial begin
			$display("B1");
	end
endmoudle
