module top;
	initial begin
			$display("B1");
		$display("B2");
	end
endmoudle
